module MEM(
    clk,
    rst_n,
    valid,
    ready,
    mode,
    in
    out
);