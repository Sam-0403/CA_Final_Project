module MY_CHIP(
    clk,
    rst_n,
    valid,
    ready,
    mode,
    in
    out
);